module instr_mem
(
    input [15:0] pc,
    output wire [31:0] instruction
);
    wire [3:0] rom_addr = pc[4:1];

    reg [15:0] rom[31:0];  
      initial  
      begin  
                rom[0] = 31'b1000000110000000;  
                rom[1] = 31'b0010110010110010;  
                rom[2] = 31'b1101110001100111;  
                rom[3] = 31'b1101110111011001;  
                rom[4] = 31'b1111110110110001;  
                rom[5] = 31'b1100000001111011; 
                rom[6] = 31'b0000000000000000;  
                rom[7] = 31'b0000000000000000;  
                rom[8] = 31'b0000000000000000;  
                rom[9] = 31'b0000000000000000;  
                rom[10] = 31'b0000000000000000;  
                rom[11] = 31'b0000000000000000;  
                rom[12] = 31'b0000000000000000;  
                rom[13] = 31'b0000000000000000;  
                rom[14] = 31'b0000000000000000;  
                rom[15] = 31'b0000000000000000;  
      end  
      assign instruction = (pc[15:0] < 32 )? rom[rom_addr[3:0]]: 16'd0;  
 endmodule   